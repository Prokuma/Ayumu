module AYUMU(
	input CLK,
	input [31:0] INPUT,
	output [31:0] OUTPUT
);

reg [10:0] CLKS;

always @(posedge CLK) begin
	case (CLKS)
		5'b00001: CLKS <= 5'b00010;
		5'b00010: CLKS <= 5'b00100;
		5'b00100: CLKS <= 5'b01000;
		5'b01000: CLKS <= 5'b10000;
		5'b10000: CLKS <= 5'b00001;
		default: CLKS <= 5'b00001;
	endcase
end

always @(posedge CLKS[2]) begin
	C_FLAG <= C_OUT;
	F_FLAG <= F_OUT;
end

initial begin
	CLKS = 4'b00001;
end

wire [15:0] NEXT;
wire [15:0] ADDR;
wire [15:0] COMMAND;

wire [3:0] CAL;
wire [1:0] MODE;
wire [7:0] IM;
wire [3:0] REG_A_ADDR;
wire [3:0] REG_B_ADDR;
wire [3:0] REG_O_ADDR;
wire [1:0] REG_O_TYPE;
wire [1:0] JUMP_MODE;
wire REG_WRITE;
wire [1:0] SEL;
wire MEM_WRITE;
wire INOUT_FLAG;

wire [127:0] REG_R;
wire [63:0] REG_IO;
wire [63:0] REG_INT;
wire [7:0] REG_A;
wire [7:0] REG_B;
wire [7:0] INT_FLAG_OUT;

reg C_FLAG;
reg F_FLAG;
wire [7:0] ALU_OUT;
wire C_OUT;
wire F_OUT;

wire [7:0] DATA;

wire INT_PROCESS;

assign OUTPUT[31:8] = REG_IO[31:8];
assign OUTPUT[7:0] = REG_IO[7:0];

PC PC(.CLK_FT(CLKS[0]), .NEXT(NEXT), .ADDR(ADDR));
ROM ROM(.ADDR(ADDR), .COMMAND(COMMAND));
DECODER DECODER(.COMMAND(COMMAND), .CAL(CAL), .MODE(MODE), .IM(IM), .REG_A(REG_A_ADDR), .REG_B(REG_B_ADDR),
															 .REG_O(REG_O_ADDR), .REG_O_TYPE(REG_O_TYPE), .JUMP_MODE(JUMP_MODE), .REG_WRITE(REG_WRITE),
															 .SEL(SEL), .MEM_WRITE(MEM_WRITE), .INOUT_FLAG(INOUT_FLAG));
REG_DC REG_DC(.CLK_DC(CLKS[1]), .REG_R(REG_R), .REG_IO(REG_IO), .SEL(SEL), .REG_O_TYPE(REG_O_TYPE), .REG_A_ADDR(REG_A_ADDR),
													.REG_B_ADDR(REG_B_ADDR), .REG_O_ADDR(REG_O_ADDR), .IM(IM), .REG_A(REG_A), .REG_B(REG_B));
ALU ALU(.CLK_EX(CLKS[2]), .IN_A(REG_A), .IN_B(REG_B), .CAL(CAL), .MODE(MODE),  .C_IN(C_FLAG), .F_IN(F_FLAG), .OUT(ALU_OUT),  .C_OUT(C_OUT), .F_OUT(F_OUT));										
MEM MEM(.CLK_MEM(CLKS[3]),  .REG_A(REG_A),.ADDR(ALU_OUT), .Q(DATA));
REG_WB REG_WB(.CLK_WB(CLKS[4]), .REG_WRITE(REG_WRITE), .F_FLAG(F_FLAG), .INOUT_FLAG(INOUT_FLAG), .INT_FLAG_OUT(INT_FLAG_OUT), .PC(ADDR), .REG_A_ADDR(REG_A_ADDR), .MODE(MODE),
													  .JUMP_MODE(JUMP_MODE), .REG_O_TYPE(REG_O_TYPE), .DATA(DATA), .INPUT(INPUT), .NEXT(NEXT), .REG_R_OUT(REG_R), .REG_IO_OUT(REG_IO), .REG_INT_FLAG_OUT(REG_INT));

INPUT_INT INPUT_0(.CLK(CLKS[4]), .INPUT(INPUT[7:0]), .INT_NO(4'd0), .REG_INT(REG_INT[7:0]), .INT_FLAG(INT_FLAG_OUT[0]));
INPUT_INT INPUT_1(.CLK(CLKS[4]), .INPUT(INPUT[15:8]), .INT_NO(4'd1), .REG_INT(REG_INT[15:8]), .INT_FLAG(INT_FLAG_OUT[1]));
INPUT_INT INPUT_2(.CLK(CLKS[4]), .INPUT(INPUT[23:16]), .INT_NO(4'd2), .REG_INT(REG_INT[23:16]), .INT_FLAG(INT_FLAG_OUT[2]));
INPUT_INT INPUT_3(.CLK(CLKS[4]), .INPUT(INPUT[31:24]), .INT_NO(4'd3), .REG_INT(REG_INT[31:24]), .INT_FLAG(INT_FLAG_OUT[3]));

TIMER_INT TIMER_0 (.CLK_WB(CLKS[4]), .REG_INT(REG_INT[39:32]),  .INT_FLAG(INT_FLAG_OUT[4]));
TIMER_INT TIMER_1 (.CLK_WB(CLKS[4]), .REG_INT(REG_INT[47:40]),  .INT_FLAG(INT_FLAG_OUT[5]));
TIMER_INT TIMER_2 (.CLK_WB(CLKS[4]), .REG_INT(REG_INT[55:48]),  .INT_FLAG(INT_FLAG_OUT[6]));
TIMER_INT TIMER_3 (.CLK_WB(CLKS[4]), .REG_INT(REG_INT[63:56]),  .INT_FLAG(INT_FLAG_OUT[7]));
													  
endmodule