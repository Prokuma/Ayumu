module ROM(
	input [15:0] ADDR,
	output reg [15:0] COMMAND
);

always @* begin
	case(ADDR)
		16'd0: COMMAND <= 16'b01011100_0000_0000;
		16'd1: COMMAND <= 16'b1000_0000_11001001;
		16'd2: COMMAND <= 16'b01100010_0100_0000;
		16'd3: COMMAND <= 16'b01011100_1000_1000;
		16'd4: COMMAND <= 16'b01011100_1100_1100;
		16'd5: COMMAND <= 16'b01011100_1101_1101;
		16'd6: COMMAND <= 16'b1000_1100_00000000;
		16'd7: COMMAND <= 16'b1000_1101_00001111;
		16'd8: COMMAND <= 16'b01010010_0100_0000;
		16'd9: COMMAND <= 16'b01000110_0000_0001;
		16'd10: COMMAND <= 16'b01011100_1100_1100;
		16'd11: COMMAND <= 16'b01011100_1101_1101;
		16'd12: COMMAND <= 16'b1000_1100_00000000;
		16'd13: COMMAND <= 16'b1000_1101_00001001;
		16'd14: COMMAND <= 16'b00010000_0000_0000;
		16'd15: COMMAND <= 16'b01000011_1000_1000;
		16'd16: COMMAND <= 16'b1000_1000_00000001;
		16'd17: COMMAND <= 16'b01000011_1100_1100;
		16'd18: COMMAND <= 16'b1000_1000_00000001;
		16'd19: COMMAND <= 16'b01000011_1101_1101;
		16'd20: COMMAND <= 16'b1000_0001_00000001;
		16'd21: COMMAND <= 16'b01000110_0000_0001;
		16'd22: COMMAND <= 16'b01000111_1101_1000;
		16'd23: COMMAND <= 16'b1001_1000_00000001;
		16'd24: COMMAND <= 16'b01000111_1100_1000;
		16'd25: COMMAND <= 16'b1001_1000_00000001;
		16'd26: COMMAND <= 16'b01000111_1000_1000;
		16'd27: COMMAND <= 16'b00010000_0010_0000;
		default: COMMAND <= 16'b01000110_0000_0001;
	 endcase
end
	
endmodule